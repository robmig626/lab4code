module state_machine_control
(
    clk,
    rst,
    start_init,
    finish_init,
    start_shuffle,
    finish_shuffle,
    write_enable_init,
    write_enable_shuffle,
    address_init,
    address_shuffle,
    
);